module simeckdecryption(inp,key,out);
input[31:0]inp;
input[15:0]key;
output[31:0]out;
wire [15:0] p1,p2,k1,k2,k3,k4,k5;

assign p2=inp[15:0];
assign p1=inp[31:16];
assign k1=(p2<<1)|(p2>>15);
assign k2=key^k1^p1;
assign k3=(p2<<5)|(p2>>11);
assign k4=p2&k3;
assign k5=k2^k4;
assign out={p2,k5};

endmodule
