module simeck32(inp,key,out);
input[31:0]inp;
input[15:0]key;
output[31:0]out;
wire [31:0] k1,k2,k3,k4,k5,k6,k7,k8,k9,k10,k11,k12,k13,k14,k15,k16,k17,k18,k19,k20,k21,k22,k23,k24,k25,k26,k27,k28,k29,k30,k31;

simeck s1(inp,key,k1);
simeck s2(k1,key,k2);
simeck s3(k2,key,k3);
simeck s4(k3,key,k4);
simeck s5(k4,key,k5);
simeck s6(k5,key,k6);
simeck s7(k6,key,k7);
simeck s8(k7,key,k8);
simeck s9(k8,key,k9);
simeck s10(k9,key,k10);
simeck s11(k10,key,k11);
simeck s12(k11,key,k12);
simeck s13(k12,key,k13);
simeck s14(k13,key,k14);
simeck s15(k14,key,k15);
simeck s16(k15,key,k16);
simeck s17(k16,key,k17);
simeck s18(k17,key,k18);
simeck s19(k18,key,k19);
simeck s20(k19,key,k20);
simeck s21(k20,key,k21);
simeck s22(k21,key,k22);
simeck s23(k22,key,k23);
simeck s24(k23,key,k24);
simeck s25(k24,key,k25);
simeck s26(k25,key,k26);
simeck s27(k26,key,k27);
simeck s28(k27,key,k28);
simeck s29(k28,key,k29);
simeck s30(k29,key,k30);
simeck s31(k30,key,k31);
simeck s32(k31,key,out);
endmodule
